/* Test of the first file 
   */

module test;

endmodule
